// megafunction wizard: %ALTSQRT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSQRT 

// ============================================================
// File Name: sqrt_int_64.v
// Megafunction Name(s):
// 			ALTSQRT
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// ************************************************************


//Copyright (C) 2020  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and any partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details, at
//https://fpgasoftware.intel.com/eula.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module sqrt_int_64 (
	aclr,
	clk,
	ena,
	radical,
	q,
	remainder);

	input	  aclr;
	input	  clk;
	input	  ena;
	input	[127:0]  radical;
	output	[63:0]  q;
	output	[64:0]  remainder;

	wire [63:0] sub_wire0;
	wire [64:0] sub_wire1;
	wire [63:0] q = sub_wire0[63:0];
	wire [64:0] remainder = sub_wire1[64:0];

	altsqrt	ALTSQRT_component (
				.aclr (aclr),
				.clk (clk),
				.ena (ena),
				.radical (radical),
				.q (sub_wire0),
				.remainder (sub_wire1));
	defparam
		ALTSQRT_component.pipeline = 2,
		ALTSQRT_component.q_port_width = 64,
		ALTSQRT_component.r_port_width = 65,
		ALTSQRT_component.width = 128;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone 10 LP"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: PIPELINE NUMERIC "2"
// Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "64"
// Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "65"
// Retrieval info: CONSTANT: WIDTH NUMERIC "128"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
// Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL "clk"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT NODEFVAL "ena"
// Retrieval info: USED_PORT: q 0 0 64 0 OUTPUT NODEFVAL "q[63..0]"
// Retrieval info: USED_PORT: radical 0 0 128 0 INPUT NODEFVAL "radical[127..0]"
// Retrieval info: USED_PORT: remainder 0 0 65 0 OUTPUT NODEFVAL "remainder[64..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @radical 0 0 128 0 radical 0 0 128 0
// Retrieval info: CONNECT: q 0 0 64 0 @q 0 0 64 0
// Retrieval info: CONNECT: remainder 0 0 65 0 @remainder 0 0 65 0
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_int_64.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_int_64.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_int_64.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_int_64.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_int_64_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_int_64_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
